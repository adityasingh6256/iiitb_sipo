
`timescale 1ns/1ps
module iiitb_sipo_tb();
reg d,clk;
wire [3:0]q;
sipo a(d, clk, q);
 
initial
begin
$dumpfile ("sipo.vcd");
 $dumpvars (0,iiitb_sipo_tb);

clk=1'b0;
forever #5 clk=~clk;
end
initial
begin
d=1;
#10 d=0;
#10 d=1;
#10 d=1;
#40 $finish;
end 
endmodule
